`timescale 1ps / 1ps

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Assume `timescale 1ps/1ps. Generate a 25 MHz square wave waveform for the Signal clk.
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module Assignment22;

logic clk = 0;

always begin
    #20000;
    clk = !clk;
end

endmodule
