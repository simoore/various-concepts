interface spi_if;
    logic clk;
    logic newd;
    logic rst;
    logic [11:0] din;
    logic sclk;
    logic cs;
    logic mosi;
endinterface